library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;
use ieee.numeric_std.all;

entity rams is
generic ( g_adress_width: integer:= 18;
          g_ram_size: integer:= 1000
        );
 port(
    clka : in std_logic;
    clkb : in std_logic;
    wea : in std_logic;
    web : in std_logic;
    addra : in std_logic_vector(g_adress_width-1 downto 0);
    addrb : in std_logic_vector(g_adress_width-1 downto 0);
    dia : in std_logic_vector(15 downto 0);
    dib : in std_logic_vector(15 downto 0);
    doa : out std_logic_vector(15 downto 0);
    dob : out std_logic_vector(15 downto 0));
end rams;
architecture syn of rams is
    type ram_type is array (g_ram_size-1 downto 0) of std_logic_vector(15 downto 0);
     signal RAM : ram_type;
   begin
 process (CLKA)
 begin
    if CLKA'event and CLKA = '1' then
            DOA <= RAM(to_integer(unsigned(ADDRA)));
            if WEA = '1' then --always 0
                    RAM(to_integer(unsigned(ADDRA))) <= DIA; --does not happen
        end if;

    end if;

    if CLKA'event and CLKA = '1' then
        DOB <= RAM(to_integer(unsigned(ADDRB)));
        if WEB = '1' then
            RAM(to_integer(unsigned(ADDRB))) <= DIB;
    end if;
 end if;

 end process;
end syn; 
